** Profile: "AC_ANALYSIS-AC_Octave"  [ d:\cadence\spb_16.6\tools\capture\tclscripts\caplearningresources\hybrid\supportfiles\analysesusingpspice\analysesusingpspice\designfiles\analysesusingpspice-PSpiceFiles\AC_ANALYSIS\AC_Octave.sim ] 

** Creating circuit file "AC_Octave.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\nitint\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 10 100k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\AC_ANALYSIS.net" 


.END
